`include "InputBuffer.sv"
`include "IsolationTreeStateMachine.sv"


module i_tree(
    input wire clk,
    input wire reset,
    input wire sensor_data, // Sensor data input to the system
    output wire anomaly_detected // Output signal indicating anomaly detection
);

// Internal connections
wire [7:0] data_from_buffer;
wire data_ready, data_processed;

// Instantiate InputBuffer
InputBuffer #(
    .DATA_WIDTH(8)
) input_buffer_inst (
    .clk(clk),
    .reset(reset),
    .sensor_data(sensor_data),
    .data_processed(data_processed), // Acknowledgment from IsolationTreeStateMachine
    .data_output(data_from_buffer),
    .data_ready(data_ready)
);

// Instantiate IsolationTreeStateMachine
IsolationTreeStateMachine isolation_tree_state_machine_inst (
    .clk(clk),
    .reset(reset),
    .data_input(data_from_buffer),
    .data_valid(data_ready),
    .anomaly_detected(anomaly_detected),
    .data_processed(data_processed) // Sends acknowledgment back to InputBuffer
);

endmodule
